`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// Company: https://shzeng.cn
// Engineer: Theo Tsang <sihao.tsang@gmail.com>
//
// Create Date: 10/09/2024 22:13:20
// Design Name: regs
// Module Name: regs
// Target Device: <target device>
// Tool versions: <tool_versions>
// Description:
//    <Description here>
// Dependencies:
//    <Dependencies here>
// Revision:
//    <Code_revision_information>
// Additional Comments:
//    <Additional_comments>
////////////////////////////////////////////////////////////////////////////////

module regs (
    // Define your module ports and parameters here
);

////////////////////////////////////////////////////////////////////
//                               main                               
////////////////////////////////////////////////////////////////////

endmodule
