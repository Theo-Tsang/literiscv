`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// Company: https://shzeng.cn
// Engineer: Theo Tsang <sihao.tsang@gmail.com>
//
// Create Date: 10/07/2024 15:17:18
// Design Name: literiscv
// Module Name: literiscv
// Target Device: <target device>
// Tool versions: <tool_versions>
// Description:
//    <Description here>
// Dependencies:
//    <Dependencies here>
// Revision:
//    <Code_revision_information>
// Additional Comments:
//    <Additional_comments>
////////////////////////////////////////////////////////////////////////////////

module literiscv (
    // Define your module ports and parameters here
);



////////////////////////////////////////////////////////////////////
//                               main                               
////////////////////////////////////////////////////////////////////





endmodule
