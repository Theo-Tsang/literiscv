`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// Company: https://shzeng.cn
// Engineer: Theo Tsang <sihao.tsang@gmail.com>
//
// Create Date: 10/09/2024 22:56:05
// Design Name: execute
// Module Name: execute
// Target Device: <target device>
// Tool versions: <tool_versions>
// Description:
//    <Description here>
// Dependencies:
//    <Dependencies here>
// Revision:
//    <Code_revision_information>
// Additional Comments:
//    <Additional_comments>
////////////////////////////////////////////////////////////////////////////////

module execute (
    // from id
    input  logic [InstDataBus - 1:              0] i_inst_data    , // instruction data, 32-bit, from id
    input  logic [InstAddrBus - 1:              0] i_inst_addr    , // instruction address, 32-bit, from id
);






endmodule
